download the latest CFME appliance for aws at access.redhat.com
